-- hazard_detection.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: Unit that detects and deals with various hazards in a
-- MIPS pipelined processor.
--
-- AUTHOR: Daniel Limanowski
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity hazard_detection is
    port(TODO);
end hazard_detection;

architecture structural of hazard_detection is

-- TODO

begin
    -- TODO

end structural;
