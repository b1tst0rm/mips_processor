-- forwarding_logic.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: Unit that processes forwarding for data hazard avoidance.
-- This unit sits in the EX (Execute) stage of a MIPS Pipelined processor.
--
-- AUTHOR: Daniel Limanowski
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity forwarding_logic is
    port(TODO);
end forwarding_logic;

architecture structural of forwarding_logic is

-- TODO

begin
    -- TODO

end structural;
